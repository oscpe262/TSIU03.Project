-- Author: Philip Johansson, Niklas Blomqvist
-- Date: October 22 2015 
-- Description: Application for analysing sound.
--	Group 41.
-- Approved by 


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity Analysis is
	port(clk,rstn		: in std_logic; 					--System signals
			lrsel 		: in std_logic; 					--Sound signal, left/right select
			LDAC,RDAC	: in signed(15 downto 0);		--Sound signal
			vsync 		: in std_logic;					--Timing signal
			lbar 			: out unsigned(7 downto 0);	--Outgoing signal to indicate how to draw the bar
			rbar			: out unsigned(7 downto 0));	--
end entity;

architecture analarch of Analysis is
	signal lrsel_old, lrsel_change 	: std_logic := '0';			--Detect new sample
	signal ildac, irdac 					: signed(15 downto 0);		--Internal signals for left/right dac
	signal lafter, rafter, temp		: unsigned(41 downto 0); 	--?? 
	signal counter							: unsigned(5 downto 0) := "101010"; -- 4
	signal vsync_old, vsync_change 	: std_logic := '0';
	
	type state_type is (s_idle, s_2, s_3);
	signal current_s: state_type := s_idle;
	
	begin
		-- Read sound signal, every 1024 clockcycle
		ildac <= LDAC;	
		irdac <= RDAC;

		process(clk, rstn) begin
			if rstn = '0' then
				lrsel_change <= '0';
				lrsel_old <= '0';
				current_s <= s_idle;
				lafter <= (others => '0');
				rafter <= (others => '0');
				temp <= (others => '0');
			elsif rising_edge(clk) then
				lrsel_old <= lrsel;			
				lrsel_change <= lrsel_old xor lrsel;
				vsync_old <= vsync;
				vsync_change <= vsync_old xor vsync;
				
				-- Detect if change has been, and if its on right or left. correct! 
				if lrsel_change = '1' and lrsel = '1' then -- Left
					lafter <= lafter - lafter(lafter'left downto 12) + unsigned(ildac * ildac);
				elsif lrsel_change = '1' and lrsel = '0' then -- Right
					rafter <= rafter - rafter(rafter'left downto 12) + unsigned(irdac * irdac);
				end if;
				
				if vsync_change = '1' and vsync = '0' then
					current_s <= s_2;
				end if;
				
				if current_s = s_idle then
					counter <= "101010";
				elsif current_s = s_2 then
					if lrsel = '1' then
						temp <= lafter;
					elsif lrsel = '0' then
						temp <= rafter;
					end if;
					
					current_s <= s_3;
				elsif current_s = s_3 then
					if temp(41) /= '1' then
						counter <= counter - 1;
						temp <= temp(40 downto 0) & "1"; 
					else
						if lrsel = '1' then
							lbar <= counter & temp(41 downto 40); 
						else
							rbar <= counter & temp(41 downto 40);
						end if;
						
						current_s <= s_idle;
					end if;
				end if;
			end if;
		end process;
end architecture;