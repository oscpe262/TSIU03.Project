library ieee;
library work;
use work.all;
use ieee.std_logic_1164.all;
-- use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

library work;

entity TB_bar_tender is
end entity;

architecture sim of TB_bar_tender is 
  COMPONENT bar_tender
 	port   (balance_input	: in signed(3 downto 0);   -- -5 to 5
			volume_input	: in unsigned(3 downto 0); -- 0 to 0
			L_bar			: in unsigned(7 downto 0); -- 0 to 171
			R_bar			: in unsigned(7 downto 0); --:--
			L_new_bar		: in unsigned(7 downto 0); --:--
			R_new_bar		: in unsigned(7 downto 0); --:--
			hcnt			: in unsigned(9 downto 0);
			vcnt			: in unsigned(9 downto 0);
			mute			: in std_logic;
			clk     		: in std_logic;
			vsync			: out std_logic;
			render_bars		: out std_logic;
			render_peak		: out std_logic;
			reset        : in  std_logic);
		end component;

	signal          balance_input : signed(3 downto 0);-- -5 to 5
	signal		volume_input: unsigned(3 downto 0); -- 0 to 0
	signal		L_bar : unsigned(7 downto 0); -- 0 to 171
	signal		R_bar : unsigned(7 downto 0); --:--
	signal		L_new_bar : unsigned(7 downto 0); --:--
	signal		R_new_bar : unsigned(7 downto 0); --:--
	signal		hcnt : unsigned(9 downto 0) := (others => '0');
	signal		vcnt : unsigned(9 downto 0) := (others => '0');
	signal		mute : std_logic;
	signal   clk : std_logic;
	signal		vsync : std_logic;
	signal		render_bars : std_logic;
	signal		render_peak : std_logic;
	signal  reset       : std_logic;

		
begin
  DUT: entity work.bar_tender port map(
  balance_input => balance_input,
  volume_input  => volume_input,
  L_bar 		=> L_bar, 
  R_bar			=> R_bar,  
  L_new_bar		=> L_new_bar,
  R_new_bar		=> R_new_bar,
  hcnt			=> hcnt, 
  vcnt			=> vcnt,
  mute			=> mute,
  clk     => clk,
  vsync			=> vsync, 
  render_bars	=> render_bars,
  render_peak	=> render_peak,
  reset => reset
  ); 
  
 balance_input <= "0101";
 volume_input <= "0101";
 L_bar <= "00000000"; --"10101010";
 R_bar <= "00000000"; --"10101010";
 L_new_bar <= "00000000"; --"10101010";
 R_new_bar <= "00000000";-- "10101010";
 mute <= '0';
 
 
 process begin
	for i in 1 to 608321 loop
	 if(clk = '0' or clk = '1') then
	   clk <= not clk;
	 else
	    clk <= '1';
	 end if;
	 
	 if(clk = '1') then
		if(hcnt < 641) then
			hcnt <= hcnt + 1;
		else 
			hcnt <= (others => '0');
		end if;
		
		if(hcnt = 640) then
		  if(vcnt < 481) then
		  	vcnt <= vcnt + 1;	
		  else 
			 vcnt <= (others => '0');
	    end if;
	   end if;
	   
	  end if;
	 wait for 50 ns;
  end loop;
end process;

	

end architecture; 
